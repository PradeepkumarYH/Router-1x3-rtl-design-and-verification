class dst_seqs_base extends uvm_sequence #(dst_xtn);
`uvm_object_utils(dst_seqs_base)
function new(string name="dst_seqs_base");
super.new(name);
endfunction
endclass
