class dst_xtn extends uvm_sequence_item;
`uvm_object_utils(dst_xtn)

function new(string name="dst_xtn");
super.new(name);
endfunction

endclass
